module opcodes
import storage

pub fn op_1001(mut app storage.App) {

	app.variables.builder.clear()
	
}